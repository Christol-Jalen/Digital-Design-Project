library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;
library gaisler;
use gaisler.misc.all;
library UNISIM;
use UNISIM.VComponents.all;

ENTITY AHB_bridge IS
  PORT(
    -- Clock and Reset -----------------
    clkm : IN std_logic;
    rstn : IN std_logic;
    -- AHB Master records --------------
    ahbmi : IN ahb_mst_in_type;
    ahbmo : OUT ahb_mst_out_type;
    -- ARM Cortex-M0 AHB-Lite signals -- 
    HADDR : IN std_logic_vector (31 downto 0); -- AHB transaction address
    HSIZE : IN std_logic_vector (2 downto 0); -- AHB size: byte, half-word or word
    HTRANS : IN std_logic_vector (1 downto 0); -- AHB transfer: non-sequential only
    HWDATA : IN std_logic_vector (31 downto 0); -- AHB write-data
    HWRITE : IN std_logic; -- AHB write control
    HRDATA : OUT std_logic_vector (31 downto 0); -- AHB read-data
    HREADY : OUT std_logic -- AHB stall signal
  );
END;

ARCHITECTURE structural OF AHB_bridge IS
  --declare a component for state_machine
  
  COMPONENT state_machine IS
    PORT(
      HADDR : IN std_logic_vector (31 downto 0);
      HSIZE : IN std_logic_vector (2 downto 0);
      HTRANS : IN std_logic_vector (1 downto 0);
      HWDATA : IN std_logic_vector (31 downto 0);
      HWRITE : IN std_logic;
      HREADY : OUT std_logic;
      dmai : OUT ahb_dma_in_type;
      dmao : IN ahb_dma_out_type; 
      clkm : IN  std_logic;
      rstn : IN std_logic
    );
  END COMPONENT;  
  
  --declare a component for ahbmstclkm
  COMPONENT ahbmst IS
    PORT(
      ahbo : OUT ahb_mst_out_type;
      ahbi : IN ahb_mst_in_type;
      dmai : IN ahb_dma_in_type;
      dmao : OUT ahb_dma_out_type;
      clk : IN  std_logic;
      rst : IN std_logic
    );
  END COMPONENT; 
  
  --declare a component for data_swapper
  COMPONENT data_swapper IS
    PORT(
      dmao : IN ahb_dma_out_type;
      HRDATA : OUT std_logic_vector (31 downto 0)
    );
  END COMPONENT; 


  SIGNAL sig_dmai : ahb_dma_in_type;
  SIGNAL sig_dmao : ahb_dma_out_type;
  SIGNAL sig_clk : std_logic;
  SIGNAL sig_rst : std_logic;
  SIGNAL sig_HADDR : std_logic_vector (31 downto 0);
  SIGNAL sig_HSIZE : std_logic_vector (2 downto 0);
  SIGNAL sig_HTRANS : std_logic_vector (1 downto 0);
  SIGNAL sig_HWDATA : std_logic_vector (31 downto 0);
  SIGNAL sig_HWRITE : std_logic;
  SIGNAL sig_HREADY : std_logic;
  SIGNAL sig_HRDATA : std_logic_vector (31 downto 0);
  SIGNAL sig_ahbo : ahb_mst_out_type;
  SIGNAL sig_ahbi : ahb_mst_in_type;


BEGIN
-----------------------------------------------------
  
  A0: ENTITY AHB_bridge
  port map(
    HADDR => sig_HADDR,
    HSIZE => sig_HSIZE,
    HTRANS => sig_HTRANS,
    HWDATA => sig_HWDATA,
    HRDATA => sig_HRDATA,
    HWRITE => sig_HWRITE,
    HREADY => sig_HREADY,
    
    ahbmi => sig_ahbi,
    ahbmo => sig_ahbo,
    
    clkm => sig_clk,
    rstn => sig_rst
  );
  
  A1: state_machine
  port map(
    HADDR => sig_HADDR,
    HSIZE => sig_HSIZE,
    HTRANS => sig_HTRANS,
    HWDATA => sig_HWDATA,
    HWRITE => sig_HWRITE,
    HREADY => sig_HREADY,
    
    dmai => sig_dmai,
    dmao => sig_dmao,
    
    clkm => sig_clk,
    rstn => sig_rst
  ); 
--instantiate state_machine component and make the connections

  A2: ahbmst
  port map(
    ahbo => sig_ahbo,
    ahbi => sig_ahbi,
    
    dmai => sig_dmai,
    dmao => sig_dmao,
    
    clk => sig_clk,
    rst => sig_rst
  );
    
--instantiate the ahbmst component and make the connections 

  A3: data_swapper
  port map(
    dmao => sig_dmao,
    HRDATA => sig_HRDATA
  );

--instantiate the data_swapper component and make the connections

END structural;
